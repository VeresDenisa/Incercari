package DB_environment_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import DB_item_pack::*;
    import DB_sequence_pack::*;
  
    import DB_agent_pack::*;
    import DB_coverage_pack::*;
   
    `include "testbench/DB/test/environment/DB_environment_config.svh"
    `include "testbench/DB/test/environment/DB_environment.svh"
  endpackage : DB_environment_pack