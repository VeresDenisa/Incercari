covergroup CM_input_covergroup (ref CM_input_item item);
    
endgroup : CM_input_covergroup