covergroup VGA_covergroup (ref VGA_output_item item);
    
endgroup : VGA_covergroup