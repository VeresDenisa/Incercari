covergroup CM_output_covergroup (ref CM_output_item item);
    
endgroup : CM_output_covergroup