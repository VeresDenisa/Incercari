package DB_item_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    `include "src/DB/test/item/DB_item.svh"
  endpackage : DB_item_pack