package VGA_sequence_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import VGA_item_pack::*;
      
    `include "testbench/CONF/test/sequence/CONF_input_sequence.svh"

    `include "testbench/VGA/test/sequence/VGA_input_sequence.svh"
  endpackage : VGA_sequence_pack