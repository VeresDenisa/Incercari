package DB_sequence_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import DB_item_pack::*;
  
    `include "src/DB/test/sequence/DB_sequence.svh"
  endpackage : DB_sequence_pack