covergroup UART_covergroup (ref UART_output_item item);
    
endgroup : UART_covergroup