package UART_item_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "testbench/CONF/test/item/CONF_item.svh"

    `include "testbench/UART/test/item/UART_input_item.svh"
    `include "testbench/UART/test/item/UART_output_item.svh"
  endpackage : UART_item_pack