covergroup LM_covergroup (ref LM_item item);
    
endgroup : LM_covergroup