package item_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    `include "testbench/DB/test/item/DB_item.svh"
  endpackage : item_pack