package VGA_item_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    `include "testbench/CONF/test/item/CONF_item.svh"
    
    `include "testbench/VGA/test/item/VGA_input_item.svh"
    `include "testbench/VGA/test/item/VGA_output_item.svh"
  endpackage : VGA_item_pack