package DB_sequence_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import DB_item_pack::*;
  
    `include "testbench/DB/test/sequence/DB_sequence.svh"
  endpackage : DB_sequence_pack