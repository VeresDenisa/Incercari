package sequence_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import item_pack::*;
  
    `include "testbench/DB/test/sequence/DB_sequence.svh"
  endpackage : sequence_pack