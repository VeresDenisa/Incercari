package CM_item_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    `include "testbench/CM/test/item/CM_input_item.svh"
    `include "testbench/CM/test/item/CM_output_item.svh"

    `include "testbench/CONF/test/item/CONF_item.svh"
  endpackage : CM_item_pack