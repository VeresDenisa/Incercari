package LM_item_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    `include "testbench/CM/test/item/CM_output_item.svh"

    `include "testbench/LM/test/item/LM_item.svh"

    `include "testbench/UART/test/item/UART_output_item.svh"
  endpackage : LM_item_pack