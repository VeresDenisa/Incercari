package CD_coverage_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import CD_item_pack::*;
  
    `include "testbench/CD/test/environment/coverage/CD_covergroup.sv"

    `include "testbench/CD/test/environment/coverage/CD_coverage.svh"
  endpackage : CD_coverage_pack