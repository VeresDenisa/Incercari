package CD_item_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    `include "testbench/CD/test/item/CD_item.svh"

    `include "testbench/CONF/test/item/CONF_item.svh"

    `include "testbench/CM/test/item/CM_input_item.svh"
  endpackage : CD_item_pack