covergroup CONF_covergroup (ref CONF_item item);
    
endgroup : CONF_covergroup